module AND_ALU (input logic [7:0] A,B, output logic [7:0] R);
    assign R = A & B;
endmodule
